module andDemo (a,b,c);

	input a,b;
	output c;

	wire a,b;
	wire c;

	assign c=a & b;

endmodule
